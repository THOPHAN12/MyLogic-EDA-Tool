module arithmetic_operations(a, b, c, d, sum_out, diff_out, prod_out, quot_out);
  input [3:0] a, b, c, d;
  output [4:0] sum_out, diff_out;
  output [7:0] prod_out;
  output [3:0] quot_out;
  
  assign sum_out = a + b;      // Addition
  assign diff_out = c - d;     // Subtraction  
  assign prod_out = a * b;     // Multiplication
  assign quot_out = c / d;     // Division
endmodule
