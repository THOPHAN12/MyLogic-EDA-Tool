/*
 * Simple AND gate test case
 * Input: a, b
 * Output: out = a & b
 */

module simple_and (
    input a,
    input b,
    output out
);

assign out = a & b;

endmodule
